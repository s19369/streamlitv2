�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.1qubX   n_estimatorsqK
X   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   objawyq0X   wiekq1X   chorobyq2X   wzrostq3etq4bX   n_features_in_q5KX
   n_outputs_q6KX   classes_q7h"h#K �q8h%�q9Rq:(KK�q;h)X   i8q<���q=Rq>(KX   <q?NNNJ����J����K tq@b�C               qAtqBbX
   n_classes_qCKX   base_estimator_qDhX   estimators_qE]qF(h)�qG}qH(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h5Kh6Kh7h"h#K �qIh%�qJRqK(KK�qLh)X   f8qM���qNRqO(Kh?NNNJ����J����K tqPb�C              �?qQtqRbhCcnumpy.core.multiarray
scalar
qSh>C       qT�qURqVX   max_features_qWKX   tree_qXcsklearn.tree._tree
Tree
qYKh"h#K �qZh%�q[Rq\(KK�q]h>�C       q^tq_bK�q`Rqa}qb(hKX
   node_countqcK	X   nodesqdh"h#K �qeh%�qfRqg(KK	�qhh)X   V56qi���qjRqk(Kh-N(X
   left_childqlX   right_childqmX   featureqnX	   thresholdqoX   impurityqpX   n_node_samplesqqX   weighted_n_node_samplesqrtqs}qt(hlh>K �quhmh>K�qvhnh>K�qwhohOK�qxhphOK �qyhqh>K(�qzhrhOK0�q{uK8KKtq|b�B�                              @     ��?             H@������������������������       �                     9@                          �E@���}<S�?             7@                            @z�G�z�?	             $@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@q}tq~bX   valuesqh"h#K �q�h%�q�Rq�(KK	KK�q�hO�C�      ;@      5@      9@               @      5@       @       @       @      �?              �?       @                      @              *@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h5Kh6Kh7h"h#K �q�h%�q�Rq�(KK�q�hO�C              �?q�tq�bhChSh>C       q��q�Rq�hWKhXhYKh"h#K �q�h%�q�Rq�(KK�q�h>�C       q�tq�bK�q�Rq�}q�(hKhcKhdh"h#K �q�h%�q�Rq�(KK�q�hk�Bh                              @�q�q��?!             H@������������������������       �        	             ,@       
                     @��hJ,�?             A@       	                    @�eP*L��?	             &@                          �@@r�q��?             @������������������������       �                     @                           C@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     7@q�tq�bhh"h#K �q�h%�q�Rq�(KKKK�q�hO�C�      3@      =@      ,@              @      =@      @      @      @      �?      @               @      �?              �?       @                      @              7@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h5Kh6Kh7h"h#K �q�h%�q�Rq�(KK�q�hO�C              �?q�tq�bhChSh>C       q��q�Rq�hWKhXhYKh"h#K �q�h%�q�Rq�(KK�q�h>�C       q�tq�bK�q�Rq�}q�(hKhcK	hdh"h#K �q�h%�q�Rq�(KK	�q�hk�B�                              @�q�q��?             H@������������������������       �                     .@                            @<���D�?            �@@                          Pf@X�<ݚ�?             "@������������������������       �                     @                           C@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@q�tq�bhh"h#K �q�h%�q�Rq�(KK	KK�q�hO�C�      3@      =@      .@              @      =@      @      @              @      @       @               @      @                      8@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h5Kh6Kh7h"h#K �q�h%�q�Rq�(KK�q�hO�C              �?q�tq�bhChSh>C       qΆq�Rq�hWKhXhYKh"h#K �q�h%�q�Rq�(KK�q�h>�C       q�tq�bK�q�Rq�}q�(hKhcKhdh"h#K �q�h%�q�Rq�(KK�q�hk�Bh                              @�q���?             H@������������������������       �                     3@       
                     @\-��p�?             =@                         ��f@�q�q�?             (@������������������������       �                     @                           C@�q�q�?             @������������������������       �                      @       	                  y
F@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     1@q�tq�bhh"h#K �q�h%�q�Rq�(KKKK�q�hO�C�      7@      9@      3@              @      9@      @       @              @      @       @       @               @       @               @       @                      1@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h5Kh6Kh7h"h#K �q�h%�q�Rq�(KK�q�hO�C              �?q�tq�bhChSh>C       q�q�Rq�hWKhXhYKh"h#K �q�h%�q�Rq�(KK�q�h>�C       q�tq�bK�q�Rq�}q�(hKhcKhdh"h#K �q�h%�q�Rq�(KK�q�hk�B�                              @�q�q�?#             H@������������������������       �                     2@                            @��S�ۿ?             >@                          �0@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@q�tq�bhh"h#K �r   h%�r  Rr  (KKKK�r  hO�Cp      4@      <@      2@               @      <@       @      @       @                      @              8@r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h5Kh6Kh7h"h#K �r  h%�r	  Rr
  (KK�r  hO�C              �?r  tr  bhChSh>C       r  �r  Rr  hWKhXhYKh"h#K �r  h%�r  Rr  (KK�r  h>�C       r  tr  bK�r  Rr  }r  (hKhcKhdh"h#K �r  h%�r  Rr  (KK�r  hk�B�                             '@     ��?             H@������������������������       �                      @                           @(옄��?             G@                            @�4�����?             ?@       
                    C@���7�?             6@                            @�����H�?             "@������������������������       �                     @       	                   �@@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             *@������������������������       �                     "@������������������������       �                     .@r  tr  bhh"h#K �r   h%�r!  Rr"  (KKKK�r#  hO�C�      5@      ;@               @      5@      9@      5@      $@      5@      �?       @      �?      @              @      �?      @                      �?      *@                      "@              .@r$  tr%  bubhhubh)�r&  }r'  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h5Kh6Kh7h"h#K �r(  h%�r)  Rr*  (KK�r+  hO�C              �?r,  tr-  bhChSh>C       r.  �r/  Rr0  hWKhXhYKh"h#K �r1  h%�r2  Rr3  (KK�r4  h>�C       r5  tr6  bK�r7  Rr8  }r9  (hKhcKhdh"h#K �r:  h%�r;  Rr<  (KK�r=  hk�BH                            �d@�q�q�?             H@������������������������       �                     @                            @���X�K�?            �F@������������������������       �                      @                          �0@$G$n��?            �B@                            @      �?             @������������������������       �                     @������������������������       �                     �?	                            @�FVQ&�?            �@@
                           @�<ݚ�?             "@                           �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     8@r>  tr?  bhh"h#K �r@  h%�rA  RrB  (KKKK�rC  hO�C�      0@      @@      @              *@      @@       @              @      @@      @      �?      @                      �?       @      ?@       @      @       @      @              @       @                      @              8@rD  trE  bubhhubh)�rF  }rG  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h5Kh6Kh7h"h#K �rH  h%�rI  RrJ  (KK�rK  hO�C              �?rL  trM  bhChSh>C       rN  �rO  RrP  hWKhXhYKh"h#K �rQ  h%�rR  RrS  (KK�rT  h>�C       rU  trV  bK�rW  RrX  }rY  (hKhcKhdh"h#K �rZ  h%�r[  Rr\  (KK�r]  hk�B�                              @      �?             H@������������������������       �                     4@                          @@@؇���X�?             <@                            @      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     4@r^  tr_  bhh"h#K �r`  h%�ra  Rrb  (KKKK�rc  hO�Cp      8@      8@      4@              @      8@      @      @      @                      @              4@rd  tre  bubhhubh)�rf  }rg  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h5Kh6Kh7h"h#K �rh  h%�ri  Rrj  (KK�rk  hO�C              �?rl  trm  bhChSh>C       rn  �ro  Rrp  hWKhXhYKh"h#K �rq  h%�rr  Rrs  (KK�rt  h>�C       ru  trv  bK�rw  Rrx  }ry  (hKhcKhdh"h#K �rz  h%�r{  Rr|  (KK�r}  hk�B�                           ��f@r�qG�?             H@                            @ҳ�wY;�?             1@������������������������       �                     &@������������������������       �                     @                            @�n`���?             ?@������������������������       �                     @                            @�>����?             ;@       	                    7@�q�q�?             @������������������������       �                     �?
                           h@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     5@r~  tr  bhh"h#K �r�  h%�r�  Rr�  (KKKK�r�  hO�C�      1@      ?@      &@      @      &@                      @      @      9@      @               @      9@       @      @      �?              �?      @              @      �?                      5@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h5Kh6Kh7h"h#K �r�  h%�r�  Rr�  (KK�r�  hO�C              �?r�  tr�  bhChSh>C       r�  �r�  Rr�  hWKhXhYKh"h#K �r�  h%�r�  Rr�  (KK�r�  h>�C       r�  tr�  bK�r�  Rr�  }r�  (hKhcKhdh"h#K �r�  h%�r�  Rr�  (KK�r�  hk�Bh                              @r�q��?             H@������������������������       �        
             3@                          �0@ܷ��?��?             =@                           '@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �h@ ��WV�?             :@������������������������       �                     3@	       
                     @؇���X�?             @������������������������       �                     �?������������������������       �                     @r�  tr�  bhh"h#K �r�  h%�r�  Rr�  (KKKK�r�  hO�C�      6@      :@      3@              @      :@       @      �?              �?       @              �?      9@              3@      �?      @      �?                      @r�  tr�  bubhhubehhub.